/escnfs/courses/sp24-cse-60762.01/public/intel16libs/pdk224_r0.9.2/apr/cadence/m11_1x_3xa_1xb_1xc_2yb_2ga_mim2_1gb__bumpp/6t108_tp0/p1222.lef