########
VERSION 5.8 ;
PROPERTYDEFINITIONS
  LIBRARY LEF58_STACKVIALAYERRULE STRING "
    STACKVIALAYERRULE via2_1x2 LAYER v2 ROWCOL 1 2 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 3 ;
    STACKVIALAYERRULE via3_2x2 LAYER v3 ROWCOL 2 2 XPITCH 2 YPITCH 2 MAXCELLEXTENSION 3 ;
    STACKVIALAYERRULE via4_2x2 LAYER v4 ROWCOL 2 1 XPITCH 1 YPITCH 1 MAXCELLEXTENSION 3 ;
  " ;

  LIBRARY LEF58_STACKVIARULE STRING "
    STACKVIARULE VP_SECPG_M1M5 via2_1x2 via3_2x2 via4_2x2 ;
  " ;
  
END PROPERTYDEFINITIONS 
############################################
