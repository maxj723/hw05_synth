/escnfs/courses/sp24-cse-60762.01/public/intel16libs/std_cells/base_nom/lef/lib224_b0m_6t_108pp_base_nom.lef