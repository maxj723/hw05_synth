/escnfs/courses/sp24-cse-60762.01/public/intel16libs/std_cells/seq_nom/lef/lib224_b0m_6t_108pp_seq_nom.lef